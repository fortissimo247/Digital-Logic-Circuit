`timescale 1ns / 1ps

module cpu_tb;

initial begin
    #20;
    $stop;
end

endmodule
